`timescale 1ns / 1ps
module tb_top();
    reg clk;
    reg reset;

    top_module dut (.clk(clk), .reset(reset));

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    initial begin
        reset = 1;
        #20;
        reset = 0;
        #800;
        $finish;
    end
endmodule
